magic
tech sky130A
magscale 1 2
timestamp 1647702129
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 14 1912 119218 117552
<< metal2 >>
rect -10 119200 102 120000
rect 2566 119200 2678 120000
rect 4498 119200 4610 120000
rect 6430 119200 6542 120000
rect 9006 119200 9118 120000
rect 10938 119200 11050 120000
rect 12870 119200 12982 120000
rect 14802 119200 14914 120000
rect 17378 119200 17490 120000
rect 19310 119200 19422 120000
rect 21242 119200 21354 120000
rect 23818 119200 23930 120000
rect 25750 119200 25862 120000
rect 27682 119200 27794 120000
rect 29614 119200 29726 120000
rect 32190 119200 32302 120000
rect 34122 119200 34234 120000
rect 36054 119200 36166 120000
rect 38630 119200 38742 120000
rect 40562 119200 40674 120000
rect 42494 119200 42606 120000
rect 45070 119200 45182 120000
rect 47002 119200 47114 120000
rect 48934 119200 49046 120000
rect 50866 119200 50978 120000
rect 53442 119200 53554 120000
rect 55374 119200 55486 120000
rect 57306 119200 57418 120000
rect 59882 119200 59994 120000
rect 61814 119200 61926 120000
rect 63746 119200 63858 120000
rect 65678 119200 65790 120000
rect 68254 119200 68366 120000
rect 70186 119200 70298 120000
rect 72118 119200 72230 120000
rect 74694 119200 74806 120000
rect 76626 119200 76738 120000
rect 78558 119200 78670 120000
rect 81134 119200 81246 120000
rect 83066 119200 83178 120000
rect 84998 119200 85110 120000
rect 86930 119200 87042 120000
rect 89506 119200 89618 120000
rect 91438 119200 91550 120000
rect 93370 119200 93482 120000
rect 95946 119200 96058 120000
rect 97878 119200 97990 120000
rect 99810 119200 99922 120000
rect 101742 119200 101854 120000
rect 104318 119200 104430 120000
rect 106250 119200 106362 120000
rect 108182 119200 108294 120000
rect 110758 119200 110870 120000
rect 112690 119200 112802 120000
rect 114622 119200 114734 120000
rect 117198 119200 117310 120000
rect 119130 119200 119242 120000
rect -10 0 102 800
rect 1922 0 2034 800
rect 3854 0 3966 800
rect 5786 0 5898 800
rect 8362 0 8474 800
rect 10294 0 10406 800
rect 12226 0 12338 800
rect 14802 0 14914 800
rect 16734 0 16846 800
rect 18666 0 18778 800
rect 20598 0 20710 800
rect 23174 0 23286 800
rect 25106 0 25218 800
rect 27038 0 27150 800
rect 29614 0 29726 800
rect 31546 0 31658 800
rect 33478 0 33590 800
rect 36054 0 36166 800
rect 37986 0 38098 800
rect 39918 0 40030 800
rect 41850 0 41962 800
rect 44426 0 44538 800
rect 46358 0 46470 800
rect 48290 0 48402 800
rect 50866 0 50978 800
rect 52798 0 52910 800
rect 54730 0 54842 800
rect 56662 0 56774 800
rect 59238 0 59350 800
rect 61170 0 61282 800
rect 63102 0 63214 800
rect 65678 0 65790 800
rect 67610 0 67722 800
rect 69542 0 69654 800
rect 72118 0 72230 800
rect 74050 0 74162 800
rect 75982 0 76094 800
rect 77914 0 78026 800
rect 80490 0 80602 800
rect 82422 0 82534 800
rect 84354 0 84466 800
rect 86930 0 87042 800
rect 88862 0 88974 800
rect 90794 0 90906 800
rect 92726 0 92838 800
rect 95302 0 95414 800
rect 97234 0 97346 800
rect 99166 0 99278 800
rect 101742 0 101854 800
rect 103674 0 103786 800
rect 105606 0 105718 800
rect 108182 0 108294 800
rect 110114 0 110226 800
rect 112046 0 112158 800
rect 113978 0 114090 800
rect 116554 0 116666 800
rect 118486 0 118598 800
<< obsm2 >>
rect 158 119144 2510 119354
rect 2734 119144 4442 119354
rect 4666 119144 6374 119354
rect 6598 119144 8950 119354
rect 9174 119144 10882 119354
rect 11106 119144 12814 119354
rect 13038 119144 14746 119354
rect 14970 119144 17322 119354
rect 17546 119144 19254 119354
rect 19478 119144 21186 119354
rect 21410 119144 23762 119354
rect 23986 119144 25694 119354
rect 25918 119144 27626 119354
rect 27850 119144 29558 119354
rect 29782 119144 32134 119354
rect 32358 119144 34066 119354
rect 34290 119144 35998 119354
rect 36222 119144 38574 119354
rect 38798 119144 40506 119354
rect 40730 119144 42438 119354
rect 42662 119144 45014 119354
rect 45238 119144 46946 119354
rect 47170 119144 48878 119354
rect 49102 119144 50810 119354
rect 51034 119144 53386 119354
rect 53610 119144 55318 119354
rect 55542 119144 57250 119354
rect 57474 119144 59826 119354
rect 60050 119144 61758 119354
rect 61982 119144 63690 119354
rect 63914 119144 65622 119354
rect 65846 119144 68198 119354
rect 68422 119144 70130 119354
rect 70354 119144 72062 119354
rect 72286 119144 74638 119354
rect 74862 119144 76570 119354
rect 76794 119144 78502 119354
rect 78726 119144 81078 119354
rect 81302 119144 83010 119354
rect 83234 119144 84942 119354
rect 85166 119144 86874 119354
rect 87098 119144 89450 119354
rect 89674 119144 91382 119354
rect 91606 119144 93314 119354
rect 93538 119144 95890 119354
rect 96114 119144 97822 119354
rect 98046 119144 99754 119354
rect 99978 119144 101686 119354
rect 101910 119144 104262 119354
rect 104486 119144 106194 119354
rect 106418 119144 108126 119354
rect 108350 119144 110702 119354
rect 110926 119144 112634 119354
rect 112858 119144 114566 119354
rect 114790 119144 117142 119354
rect 117366 119144 119074 119354
rect 20 856 119212 119144
rect 158 31 1866 856
rect 2090 31 3798 856
rect 4022 31 5730 856
rect 5954 31 8306 856
rect 8530 31 10238 856
rect 10462 31 12170 856
rect 12394 31 14746 856
rect 14970 31 16678 856
rect 16902 31 18610 856
rect 18834 31 20542 856
rect 20766 31 23118 856
rect 23342 31 25050 856
rect 25274 31 26982 856
rect 27206 31 29558 856
rect 29782 31 31490 856
rect 31714 31 33422 856
rect 33646 31 35998 856
rect 36222 31 37930 856
rect 38154 31 39862 856
rect 40086 31 41794 856
rect 42018 31 44370 856
rect 44594 31 46302 856
rect 46526 31 48234 856
rect 48458 31 50810 856
rect 51034 31 52742 856
rect 52966 31 54674 856
rect 54898 31 56606 856
rect 56830 31 59182 856
rect 59406 31 61114 856
rect 61338 31 63046 856
rect 63270 31 65622 856
rect 65846 31 67554 856
rect 67778 31 69486 856
rect 69710 31 72062 856
rect 72286 31 73994 856
rect 74218 31 75926 856
rect 76150 31 77858 856
rect 78082 31 80434 856
rect 80658 31 82366 856
rect 82590 31 84298 856
rect 84522 31 86874 856
rect 87098 31 88806 856
rect 89030 31 90738 856
rect 90962 31 92670 856
rect 92894 31 95246 856
rect 95470 31 97178 856
rect 97402 31 99110 856
rect 99334 31 101686 856
rect 101910 31 103618 856
rect 103842 31 105550 856
rect 105774 31 108126 856
rect 108350 31 110058 856
rect 110282 31 111990 856
rect 112214 31 113922 856
rect 114146 31 116498 856
rect 116722 31 118430 856
rect 118654 31 119212 856
<< metal3 >>
rect 119200 118948 120000 119188
rect 0 118268 800 118508
rect 119200 116908 120000 117148
rect 0 116228 800 116468
rect 119200 114188 120000 114428
rect 0 113508 800 113748
rect 119200 112148 120000 112388
rect 0 111468 800 111708
rect 119200 110108 120000 110348
rect 0 109428 800 109668
rect 0 107388 800 107628
rect 119200 107388 120000 107628
rect 119200 105348 120000 105588
rect 0 104668 800 104908
rect 119200 103308 120000 103548
rect 0 102628 800 102868
rect 119200 101268 120000 101508
rect 0 100588 800 100828
rect 119200 98548 120000 98788
rect 0 97868 800 98108
rect 119200 96508 120000 96748
rect 0 95828 800 96068
rect 119200 94468 120000 94708
rect 0 93788 800 94028
rect 0 91748 800 91988
rect 119200 91748 120000 91988
rect 119200 89708 120000 89948
rect 0 89028 800 89268
rect 119200 87668 120000 87908
rect 0 86988 800 87228
rect 0 84948 800 85188
rect 119200 84948 120000 85188
rect 119200 82908 120000 83148
rect 0 82228 800 82468
rect 119200 80868 120000 81108
rect 0 80188 800 80428
rect 119200 78828 120000 79068
rect 0 78148 800 78388
rect 119200 76108 120000 76348
rect 0 75428 800 75668
rect 119200 74068 120000 74308
rect 0 73388 800 73628
rect 119200 72028 120000 72268
rect 0 71348 800 71588
rect 0 69308 800 69548
rect 119200 69308 120000 69548
rect 119200 67268 120000 67508
rect 0 66588 800 66828
rect 119200 65228 120000 65468
rect 0 64548 800 64788
rect 119200 63188 120000 63428
rect 0 62508 800 62748
rect 119200 60468 120000 60708
rect 0 59788 800 60028
rect 119200 58428 120000 58668
rect 0 57748 800 57988
rect 119200 56388 120000 56628
rect 0 55708 800 55948
rect 0 53668 800 53908
rect 119200 53668 120000 53908
rect 119200 51628 120000 51868
rect 0 50948 800 51188
rect 119200 49588 120000 49828
rect 0 48908 800 49148
rect 0 46868 800 47108
rect 119200 46868 120000 47108
rect 119200 44828 120000 45068
rect 0 44148 800 44388
rect 119200 42788 120000 43028
rect 0 42108 800 42348
rect 119200 40748 120000 40988
rect 0 40068 800 40308
rect 119200 38028 120000 38268
rect 0 37348 800 37588
rect 119200 35988 120000 36228
rect 0 35308 800 35548
rect 119200 33948 120000 34188
rect 0 33268 800 33508
rect 0 31228 800 31468
rect 119200 31228 120000 31468
rect 119200 29188 120000 29428
rect 0 28508 800 28748
rect 119200 27148 120000 27388
rect 0 26468 800 26708
rect 119200 25108 120000 25348
rect 0 24428 800 24668
rect 119200 22388 120000 22628
rect 0 21708 800 21948
rect 119200 20348 120000 20588
rect 0 19668 800 19908
rect 119200 18308 120000 18548
rect 0 17628 800 17868
rect 0 15588 800 15828
rect 119200 15588 120000 15828
rect 119200 13548 120000 13788
rect 0 12868 800 13108
rect 119200 11508 120000 11748
rect 0 10828 800 11068
rect 0 8788 800 9028
rect 119200 8788 120000 9028
rect 119200 6748 120000 6988
rect 0 6068 800 6308
rect 119200 4708 120000 4948
rect 0 4028 800 4268
rect 119200 2668 120000 2908
rect 0 1988 800 2228
rect 119200 -52 120000 188
<< obsm3 >>
rect 800 118868 119120 119101
rect 800 118588 119200 118868
rect 880 118188 119200 118588
rect 800 117228 119200 118188
rect 800 116828 119120 117228
rect 800 116548 119200 116828
rect 880 116148 119200 116548
rect 800 114508 119200 116148
rect 800 114108 119120 114508
rect 800 113828 119200 114108
rect 880 113428 119200 113828
rect 800 112468 119200 113428
rect 800 112068 119120 112468
rect 800 111788 119200 112068
rect 880 111388 119200 111788
rect 800 110428 119200 111388
rect 800 110028 119120 110428
rect 800 109748 119200 110028
rect 880 109348 119200 109748
rect 800 107708 119200 109348
rect 880 107308 119120 107708
rect 800 105668 119200 107308
rect 800 105268 119120 105668
rect 800 104988 119200 105268
rect 880 104588 119200 104988
rect 800 103628 119200 104588
rect 800 103228 119120 103628
rect 800 102948 119200 103228
rect 880 102548 119200 102948
rect 800 101588 119200 102548
rect 800 101188 119120 101588
rect 800 100908 119200 101188
rect 880 100508 119200 100908
rect 800 98868 119200 100508
rect 800 98468 119120 98868
rect 800 98188 119200 98468
rect 880 97788 119200 98188
rect 800 96828 119200 97788
rect 800 96428 119120 96828
rect 800 96148 119200 96428
rect 880 95748 119200 96148
rect 800 94788 119200 95748
rect 800 94388 119120 94788
rect 800 94108 119200 94388
rect 880 93708 119200 94108
rect 800 92068 119200 93708
rect 880 91668 119120 92068
rect 800 90028 119200 91668
rect 800 89628 119120 90028
rect 800 89348 119200 89628
rect 880 88948 119200 89348
rect 800 87988 119200 88948
rect 800 87588 119120 87988
rect 800 87308 119200 87588
rect 880 86908 119200 87308
rect 800 85268 119200 86908
rect 880 84868 119120 85268
rect 800 83228 119200 84868
rect 800 82828 119120 83228
rect 800 82548 119200 82828
rect 880 82148 119200 82548
rect 800 81188 119200 82148
rect 800 80788 119120 81188
rect 800 80508 119200 80788
rect 880 80108 119200 80508
rect 800 79148 119200 80108
rect 800 78748 119120 79148
rect 800 78468 119200 78748
rect 880 78068 119200 78468
rect 800 76428 119200 78068
rect 800 76028 119120 76428
rect 800 75748 119200 76028
rect 880 75348 119200 75748
rect 800 74388 119200 75348
rect 800 73988 119120 74388
rect 800 73708 119200 73988
rect 880 73308 119200 73708
rect 800 72348 119200 73308
rect 800 71948 119120 72348
rect 800 71668 119200 71948
rect 880 71268 119200 71668
rect 800 69628 119200 71268
rect 880 69228 119120 69628
rect 800 67588 119200 69228
rect 800 67188 119120 67588
rect 800 66908 119200 67188
rect 880 66508 119200 66908
rect 800 65548 119200 66508
rect 800 65148 119120 65548
rect 800 64868 119200 65148
rect 880 64468 119200 64868
rect 800 63508 119200 64468
rect 800 63108 119120 63508
rect 800 62828 119200 63108
rect 880 62428 119200 62828
rect 800 60788 119200 62428
rect 800 60388 119120 60788
rect 800 60108 119200 60388
rect 880 59708 119200 60108
rect 800 58748 119200 59708
rect 800 58348 119120 58748
rect 800 58068 119200 58348
rect 880 57668 119200 58068
rect 800 56708 119200 57668
rect 800 56308 119120 56708
rect 800 56028 119200 56308
rect 880 55628 119200 56028
rect 800 53988 119200 55628
rect 880 53588 119120 53988
rect 800 51948 119200 53588
rect 800 51548 119120 51948
rect 800 51268 119200 51548
rect 880 50868 119200 51268
rect 800 49908 119200 50868
rect 800 49508 119120 49908
rect 800 49228 119200 49508
rect 880 48828 119200 49228
rect 800 47188 119200 48828
rect 880 46788 119120 47188
rect 800 45148 119200 46788
rect 800 44748 119120 45148
rect 800 44468 119200 44748
rect 880 44068 119200 44468
rect 800 43108 119200 44068
rect 800 42708 119120 43108
rect 800 42428 119200 42708
rect 880 42028 119200 42428
rect 800 41068 119200 42028
rect 800 40668 119120 41068
rect 800 40388 119200 40668
rect 880 39988 119200 40388
rect 800 38348 119200 39988
rect 800 37948 119120 38348
rect 800 37668 119200 37948
rect 880 37268 119200 37668
rect 800 36308 119200 37268
rect 800 35908 119120 36308
rect 800 35628 119200 35908
rect 880 35228 119200 35628
rect 800 34268 119200 35228
rect 800 33868 119120 34268
rect 800 33588 119200 33868
rect 880 33188 119200 33588
rect 800 31548 119200 33188
rect 880 31148 119120 31548
rect 800 29508 119200 31148
rect 800 29108 119120 29508
rect 800 28828 119200 29108
rect 880 28428 119200 28828
rect 800 27468 119200 28428
rect 800 27068 119120 27468
rect 800 26788 119200 27068
rect 880 26388 119200 26788
rect 800 25428 119200 26388
rect 800 25028 119120 25428
rect 800 24748 119200 25028
rect 880 24348 119200 24748
rect 800 22708 119200 24348
rect 800 22308 119120 22708
rect 800 22028 119200 22308
rect 880 21628 119200 22028
rect 800 20668 119200 21628
rect 800 20268 119120 20668
rect 800 19988 119200 20268
rect 880 19588 119200 19988
rect 800 18628 119200 19588
rect 800 18228 119120 18628
rect 800 17948 119200 18228
rect 880 17548 119200 17948
rect 800 15908 119200 17548
rect 880 15508 119120 15908
rect 800 13868 119200 15508
rect 800 13468 119120 13868
rect 800 13188 119200 13468
rect 880 12788 119200 13188
rect 800 11828 119200 12788
rect 800 11428 119120 11828
rect 800 11148 119200 11428
rect 880 10748 119200 11148
rect 800 9108 119200 10748
rect 880 8708 119120 9108
rect 800 7068 119200 8708
rect 800 6668 119120 7068
rect 800 6388 119200 6668
rect 880 5988 119200 6388
rect 800 5028 119200 5988
rect 800 4628 119120 5028
rect 800 4348 119200 4628
rect 880 3948 119200 4348
rect 800 2988 119200 3948
rect 800 2588 119120 2988
rect 800 2308 119200 2588
rect 880 1908 119200 2308
rect 800 268 119200 1908
rect 800 35 119120 268
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 18091 3299 19488 95301
rect 19968 3299 34848 95301
rect 35328 3299 50208 95301
rect 50688 3299 65568 95301
rect 66048 3299 80928 95301
rect 81408 3299 96288 95301
rect 96768 3299 102797 95301
<< labels >>
rlabel metal2 s -10 119200 102 120000 6 active
port 1 nsew signal input
rlabel metal3 s 119200 35988 120000 36228 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 88862 0 88974 800 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 92726 0 92838 800 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 119200 18308 120000 18548 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 119200 13548 120000 13788 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 119200 60468 120000 60708 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 119200 44828 120000 45068 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 97234 0 97346 800 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 38630 119200 38742 120000 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 119200 2668 120000 2908 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 119200 87668 120000 87908 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 17378 119200 17490 120000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 101742 119200 101854 120000 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 0 82228 800 82468 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 110758 119200 110870 120000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 57306 119200 57418 120000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 90794 0 90906 800 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 77914 0 78026 800 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 23818 119200 23930 120000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 4498 119200 4610 120000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 32190 119200 32302 120000 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 119200 4708 120000 4948 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 63102 0 63214 800 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 119200 40748 120000 40988 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 0 109428 800 109668 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 119200 80868 120000 81108 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 101742 0 101854 800 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 0 97868 800 98108 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 52798 0 52910 800 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 99166 0 99278 800 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 80490 0 80602 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal2 s 86930 119200 87042 120000 6 io_oeb[10]
port 41 nsew signal output
rlabel metal2 s 105606 0 105718 800 6 io_oeb[11]
port 42 nsew signal output
rlabel metal2 s 91438 119200 91550 120000 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 119200 72028 120000 72268 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 119200 96508 120000 96748 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 119200 69308 120000 69548 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 0 40068 800 40308 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 59238 0 59350 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 108182 119200 108294 120000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 0 21708 800 21948 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 119200 6748 120000 6988 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 0 1988 800 2228 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 33478 0 33590 800 6 io_oeb[21]
port 53 nsew signal output
rlabel metal3 s 119200 110108 120000 110348 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 97878 119200 97990 120000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 10294 0 10406 800 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 37986 0 38098 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 119200 67268 120000 67508 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 75982 0 76094 800 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 0 37348 800 37588 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 55374 119200 55486 120000 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 0 89028 800 89268 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 10938 119200 11050 120000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 117198 119200 117310 120000 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 68254 119200 68366 120000 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 119200 103308 120000 103548 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 119200 105348 120000 105588 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 59788 800 60028 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 99810 119200 99922 120000 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 119200 76108 120000 76348 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 21242 119200 21354 120000 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 119200 33948 120000 34188 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 100588 800 100828 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 12870 119200 12982 120000 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 119200 112148 120000 112388 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 119200 58428 120000 58668 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 0 50948 800 51188 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 0 113508 800 113748 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 0 4028 800 4268 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 65678 0 65790 800 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 53668 800 53908 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 74694 119200 74806 120000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 119130 119200 119242 120000 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 80188 800 80428 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 12226 0 12338 800 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 45070 119200 45182 120000 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 119200 27148 120000 27388 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 104318 119200 104430 120000 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 0 6068 800 6308 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 0 44148 800 44388 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 103674 0 103786 800 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 114622 119200 114734 120000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 81134 119200 81246 120000 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 119200 74068 120000 74308 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 0 91748 800 91988 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 118486 0 118598 800 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 119200 51628 120000 51868 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 72118 119200 72230 120000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 89506 119200 89618 120000 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 119200 38028 120000 38268 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 8788 800 9028 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 78558 119200 78670 120000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 29614 119200 29726 120000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 48934 119200 49046 120000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 65678 119200 65790 120000 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 116554 0 116666 800 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 0 26468 800 26708 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 119200 8788 120000 9028 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 0 66588 800 66828 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 63746 119200 63858 120000 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 119200 53668 120000 53908 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 119200 22388 120000 22628 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 0 116228 800 116468 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 119200 101268 120000 101508 6 io_out[9]
port 115 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 116 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 116 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 116 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 116 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 117 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 117 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 117 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 117 nsew ground input
rlabel metal2 s 40562 119200 40674 120000 6 wb_clk_i
port 118 nsew signal input
rlabel metal3 s 119200 116908 120000 117148 6 wb_rst_i
port 119 nsew signal input
rlabel metal3 s 0 86988 800 87228 6 wbs_ack_o
port 120 nsew signal output
rlabel metal3 s 119200 78828 120000 79068 6 wbs_adr_i[0]
port 121 nsew signal input
rlabel metal3 s 119200 98548 120000 98788 6 wbs_adr_i[10]
port 122 nsew signal input
rlabel metal3 s 0 71348 800 71588 6 wbs_adr_i[11]
port 123 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 wbs_adr_i[12]
port 124 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 wbs_adr_i[13]
port 125 nsew signal input
rlabel metal3 s 119200 29188 120000 29428 6 wbs_adr_i[14]
port 126 nsew signal input
rlabel metal2 s 61814 119200 61926 120000 6 wbs_adr_i[15]
port 127 nsew signal input
rlabel metal2 s 54730 0 54842 800 6 wbs_adr_i[16]
port 128 nsew signal input
rlabel metal3 s 119200 20348 120000 20588 6 wbs_adr_i[17]
port 129 nsew signal input
rlabel metal2 s 113978 0 114090 800 6 wbs_adr_i[18]
port 130 nsew signal input
rlabel metal3 s 0 107388 800 107628 6 wbs_adr_i[19]
port 131 nsew signal input
rlabel metal3 s 0 78148 800 78388 6 wbs_adr_i[1]
port 132 nsew signal input
rlabel metal3 s 119200 65228 120000 65468 6 wbs_adr_i[20]
port 133 nsew signal input
rlabel metal3 s 0 95828 800 96068 6 wbs_adr_i[21]
port 134 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 wbs_adr_i[22]
port 135 nsew signal input
rlabel metal2 s 110114 0 110226 800 6 wbs_adr_i[23]
port 136 nsew signal input
rlabel metal2 s 36054 119200 36166 120000 6 wbs_adr_i[24]
port 137 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 wbs_adr_i[25]
port 138 nsew signal input
rlabel metal3 s 0 57748 800 57988 6 wbs_adr_i[26]
port 139 nsew signal input
rlabel metal3 s 0 75428 800 75668 6 wbs_adr_i[27]
port 140 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 wbs_adr_i[28]
port 141 nsew signal input
rlabel metal2 s 34122 119200 34234 120000 6 wbs_adr_i[29]
port 142 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 wbs_adr_i[2]
port 143 nsew signal input
rlabel metal2 s 14802 119200 14914 120000 6 wbs_adr_i[30]
port 144 nsew signal input
rlabel metal3 s 119200 11508 120000 11748 6 wbs_adr_i[31]
port 145 nsew signal input
rlabel metal2 s 72118 0 72230 800 6 wbs_adr_i[3]
port 146 nsew signal input
rlabel metal3 s 119200 94468 120000 94708 6 wbs_adr_i[4]
port 147 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 wbs_adr_i[5]
port 148 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 wbs_adr_i[6]
port 149 nsew signal input
rlabel metal2 s 25750 119200 25862 120000 6 wbs_adr_i[7]
port 150 nsew signal input
rlabel metal2 s 95302 0 95414 800 6 wbs_adr_i[8]
port 151 nsew signal input
rlabel metal3 s 0 73388 800 73628 6 wbs_adr_i[9]
port 152 nsew signal input
rlabel metal2 s 95946 119200 96058 120000 6 wbs_cyc_i
port 153 nsew signal input
rlabel metal2 s 2566 119200 2678 120000 6 wbs_dat_i[0]
port 154 nsew signal input
rlabel metal2 s 27682 119200 27794 120000 6 wbs_dat_i[10]
port 155 nsew signal input
rlabel metal2 s 47002 119200 47114 120000 6 wbs_dat_i[11]
port 156 nsew signal input
rlabel metal2 s 42494 119200 42606 120000 6 wbs_dat_i[12]
port 157 nsew signal input
rlabel metal2 s 3854 0 3966 800 6 wbs_dat_i[13]
port 158 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 wbs_dat_i[14]
port 159 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 wbs_dat_i[15]
port 160 nsew signal input
rlabel metal2 s 56662 0 56774 800 6 wbs_dat_i[16]
port 161 nsew signal input
rlabel metal3 s 119200 114188 120000 114428 6 wbs_dat_i[17]
port 162 nsew signal input
rlabel metal2 s 6430 119200 6542 120000 6 wbs_dat_i[18]
port 163 nsew signal input
rlabel metal2 s 59882 119200 59994 120000 6 wbs_dat_i[19]
port 164 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 wbs_dat_i[1]
port 165 nsew signal input
rlabel metal3 s 119200 42788 120000 43028 6 wbs_dat_i[20]
port 166 nsew signal input
rlabel metal3 s 119200 89708 120000 89948 6 wbs_dat_i[21]
port 167 nsew signal input
rlabel metal3 s 0 55708 800 55948 6 wbs_dat_i[22]
port 168 nsew signal input
rlabel metal3 s 119200 63188 120000 63428 6 wbs_dat_i[23]
port 169 nsew signal input
rlabel metal3 s 0 104668 800 104908 6 wbs_dat_i[24]
port 170 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 wbs_dat_i[25]
port 171 nsew signal input
rlabel metal3 s 119200 107388 120000 107628 6 wbs_dat_i[26]
port 172 nsew signal input
rlabel metal2 s 70186 119200 70298 120000 6 wbs_dat_i[27]
port 173 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 wbs_dat_i[28]
port 174 nsew signal input
rlabel metal3 s 119200 46868 120000 47108 6 wbs_dat_i[29]
port 175 nsew signal input
rlabel metal2 s 84354 0 84466 800 6 wbs_dat_i[2]
port 176 nsew signal input
rlabel metal3 s 119200 15588 120000 15828 6 wbs_dat_i[30]
port 177 nsew signal input
rlabel metal3 s 0 111468 800 111708 6 wbs_dat_i[31]
port 178 nsew signal input
rlabel metal2 s 108182 0 108294 800 6 wbs_dat_i[3]
port 179 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 wbs_dat_i[4]
port 180 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 wbs_dat_i[5]
port 181 nsew signal input
rlabel metal3 s 119200 31228 120000 31468 6 wbs_dat_i[6]
port 182 nsew signal input
rlabel metal3 s 119200 118948 120000 119188 6 wbs_dat_i[7]
port 183 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 wbs_dat_i[8]
port 184 nsew signal input
rlabel metal2 s 112046 0 112158 800 6 wbs_dat_i[9]
port 185 nsew signal input
rlabel metal3 s 0 46868 800 47108 6 wbs_dat_o[0]
port 186 nsew signal output
rlabel metal3 s 119200 49588 120000 49828 6 wbs_dat_o[10]
port 187 nsew signal output
rlabel metal2 s 1922 0 2034 800 6 wbs_dat_o[11]
port 188 nsew signal output
rlabel metal3 s 119200 91748 120000 91988 6 wbs_dat_o[12]
port 189 nsew signal output
rlabel metal2 s 112690 119200 112802 120000 6 wbs_dat_o[13]
port 190 nsew signal output
rlabel metal3 s 119200 -52 120000 188 6 wbs_dat_o[14]
port 191 nsew signal output
rlabel metal2 s 106250 119200 106362 120000 6 wbs_dat_o[15]
port 192 nsew signal output
rlabel metal3 s 0 64548 800 64788 6 wbs_dat_o[16]
port 193 nsew signal output
rlabel metal3 s 0 69308 800 69548 6 wbs_dat_o[17]
port 194 nsew signal output
rlabel metal2 s 74050 0 74162 800 6 wbs_dat_o[18]
port 195 nsew signal output
rlabel metal2 s -10 0 102 800 6 wbs_dat_o[19]
port 196 nsew signal output
rlabel metal2 s 86930 0 87042 800 6 wbs_dat_o[1]
port 197 nsew signal output
rlabel metal3 s 0 84948 800 85188 6 wbs_dat_o[20]
port 198 nsew signal output
rlabel metal2 s 9006 119200 9118 120000 6 wbs_dat_o[21]
port 199 nsew signal output
rlabel metal2 s 53442 119200 53554 120000 6 wbs_dat_o[22]
port 200 nsew signal output
rlabel metal3 s 0 62508 800 62748 6 wbs_dat_o[23]
port 201 nsew signal output
rlabel metal2 s 23174 0 23286 800 6 wbs_dat_o[24]
port 202 nsew signal output
rlabel metal2 s 8362 0 8474 800 6 wbs_dat_o[25]
port 203 nsew signal output
rlabel metal2 s 76626 119200 76738 120000 6 wbs_dat_o[26]
port 204 nsew signal output
rlabel metal2 s 50866 119200 50978 120000 6 wbs_dat_o[27]
port 205 nsew signal output
rlabel metal2 s 61170 0 61282 800 6 wbs_dat_o[28]
port 206 nsew signal output
rlabel metal2 s 93370 119200 93482 120000 6 wbs_dat_o[29]
port 207 nsew signal output
rlabel metal3 s 119200 25108 120000 25348 6 wbs_dat_o[2]
port 208 nsew signal output
rlabel metal3 s 0 93788 800 94028 6 wbs_dat_o[30]
port 209 nsew signal output
rlabel metal3 s 119200 84948 120000 85188 6 wbs_dat_o[31]
port 210 nsew signal output
rlabel metal2 s 25106 0 25218 800 6 wbs_dat_o[3]
port 211 nsew signal output
rlabel metal2 s 41850 0 41962 800 6 wbs_dat_o[4]
port 212 nsew signal output
rlabel metal2 s 67610 0 67722 800 6 wbs_dat_o[5]
port 213 nsew signal output
rlabel metal3 s 119200 82908 120000 83148 6 wbs_dat_o[6]
port 214 nsew signal output
rlabel metal2 s 69542 0 69654 800 6 wbs_dat_o[7]
port 215 nsew signal output
rlabel metal2 s 84998 119200 85110 120000 6 wbs_dat_o[8]
port 216 nsew signal output
rlabel metal2 s 83066 119200 83178 120000 6 wbs_dat_o[9]
port 217 nsew signal output
rlabel metal3 s 0 118268 800 118508 6 wbs_sel_i[0]
port 218 nsew signal input
rlabel metal2 s 19310 119200 19422 120000 6 wbs_sel_i[1]
port 219 nsew signal input
rlabel metal2 s 82422 0 82534 800 6 wbs_sel_i[2]
port 220 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 wbs_sel_i[3]
port 221 nsew signal input
rlabel metal3 s 0 102628 800 102868 6 wbs_stb_i
port 222 nsew signal input
rlabel metal3 s 119200 56388 120000 56628 6 wbs_we_i
port 223 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27084470
string GDS_FILE /openlane/designs/wrapped_teras/runs/RUN_2022.03.19_14.55.39/results/finishing/wrapped_teras.magic.gds
string GDS_START 1143280
<< end >>

